interface dut_if
    // declare ports here
    logic clock, reset;
    logic[7:0] portA, portB;
endinterface
