interface dut_if
    // declare ports here
endinterface
