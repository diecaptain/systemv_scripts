interface dut_if
    // declare ports here
    // logic port
    // logic [n:0] port
endinterface
